// Example 1
    #100;
    player_x = 100;
    player_y = 200;
    #100;

    // Example 2
    player_x = 50;
    player_y = 150;
    #100;

    // Example 3
    player_x = 200;
    player_y = 300;
    #100;

    // Example 4
    player_x = 80;
    player_y = 250;
    #100;

    // Example 5
    player_x = 120;
    player_y = 180;
    #100;

    // Example 6
    player_x = 60;
    player_y = 220;
    #100;

    // Example 7
    player_x = 180;
    player_y = 280;
    #100;

    // Example 8
    player_x = 90;
    player_y = 190;
    #100;

    // Example 9
    player_x = 110;
    player_y = 210;
    #100;

    // Example 10
    player_x = 70;
    player_y = 240;
    #100;

    // End simulation
    #100 $finish;
end

endmodule
